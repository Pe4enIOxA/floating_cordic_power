---------------------------------------------------------------------------
-- This VHDL file was developed by Daniel Llamocca (2013).  It may be
-- freely copied and/or distributed at no cost.  Any persons using this
-- file for any purpose do so at their own risk, and are responsible for
-- the results of such use.  Daniel Llamocca does not guarantee that
-- this file is complete, correct, or fit for any particular purpose.
-- NO WARRANTY OF ANY KIND IS EXPRESSED OR IMPLIED.  This notice must
-- accompany any copy of this file.
--------------------------------------------------------------------------
-- General N-bit Register Kazumi Malhan Final Project

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- N-bit Register
entity my_rege is
   generic (N: INTEGER:= 4);
	port ( clock, resetn: in std_logic;
	       E: in std_logic;
		  D: in std_logic_vector (N-1 downto 0);
	       Q: out std_logic_vector (N-1 downto 0));
end my_rege;

architecture Behavioral of my_rege is

	signal Qt: std_logic_vector (N-1 downto 0);
	
begin

	process (resetn, clock, E)
	begin
		if resetn = '0' then
			Qt <= (others => '0');
		elsif (clock'event and clock = '1') then
			if E = '1' then	
					Qt <= D;
			end if;
		end if;
	end process;

	Q <= Qt;
end Behavioral;

