-- LUT for npos, Kazumi Malhan, Final Project 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- LUT using multiplexer.
entity my_posLUT is
   generic (N: INTEGER:= 16);
	port (s: in std_logic_vector (3 downto 0);
	      y: out std_logic_vector (N-1 downto 0));
end my_posLUT;

architecture structure of my_posLUT is

signal a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15: std_logic_vector(N-1 downto 0);

begin
    -- These values are pre-calculated using MATLAB
bit32: if (N = 32) generate
    a0 <= x"3f0c9f54";
    a1 <= x"3e82c578";
    a2 <= x"3e00ac49";
    a3 <= x"3d802ac4";
    a4 <= x"3d000aac";
    a5 <= x"3c8002ab";
    a6 <= x"3c0000ab";
    a7 <= x"3b80002b";
    a8 <= x"3b00000b";
    a9 <= x"3a800003";
    a10 <= x"3a000001";
    a11 <= x"39800000";
    a12 <= x"39000000";
    a13 <= x"38800000";
    a14 <= x"38000000";
    a15 <= x"37800000";
    end generate;
    
bit64: if (N = 64) generate
    a0 <= x"3fe193ea7aad030b";
    a1 <= x"3fd058aefa811452";
    a2 <= x"3fc015891c9eaef7";
    a3 <= x"3fb005588ad375ad";
    a4 <= x"3fa001558891aee3";
    a5 <= x"3f9000555888ad1d";
    a6 <= x"3f8000155588891b";
    a7 <= x"3f7000055558888b";
    a8 <= x"3f60000155558889";
    a9 <= x"3f50000055555889";
    a10 <= x"3f40000015555589";
    a11 <= x"3f30000005555559";
    a12 <= x"3f20000001555556";
    a13 <= x"3f10000000555555";
    a14 <= x"3f00000000155555";
    a15 <= x"3ef0000000055555";
    end generate;
    
bit24: if (N = 24) generate
    a0 <= "001111100001100100111110";
    a1 <= "001111010000010110001010";
    a2 <= "001111000000000101011000";
    a3 <= "001110110000000001010101";
    a4 <= "001110100000000000010101";
    a5 <= "001110010000000000000101";
    a6 <= "001110000000000000000001";
    a7 <= "001101110000000000000000";
    a8 <= "001101100000000000000000";
    a9 <= "001101010000000000000000";
    a10 <= "001101000000000000000000";
    a11 <= "001100110000000000000000";
    a12 <= "001100100000000000000000";
    a13 <= "001100010000000000000000";
    a14 <= "001100000000000000000000";
    a15 <= "001011110000000000000000";
    end generate;
    
bit16: if (N = 24) generate
    a0 <= "0011110000110010";
    a1 <= "0011101000001011";
    a2 <= "0011100000000010";
    a3 <= "0011011000000000";
    a4 <= "0011010000000000";
    a5 <= "0011001000000000";
    a6 <= "0011000000000000";
    a7 <= "0010111000000000";
    a8 <= "0010111000000000";
    a9 <= "0010111000000000";
    a10 <= "0010111000000000";
    a11 <= "0010111000000000";
    a12 <= "0010111000000000";
    a13 <= "0010111000000000";
    a14 <= "0010111000000000";
    a15 <= "0010111000000000";
    end generate;
    
	with s select
		y <=   a0 when "0001",
			   a1 when "0010",
			   a2 when "0011",
			   a3 when "0100",
			   a4 when "0101",
			   a5 when "0110",
			   a6 when "0111",
			   a7 when "1000",
			   a8 when "1001",
			   a9 when "1010",
			   a10 when "1011",
			   a11 when "1100",
			   a12 when "1101",
			   a13 when "1110",
			   a14 when "1111",
			   a15 when others;
			 
end structure;